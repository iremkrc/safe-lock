----------------------------------------------------------------------------------
-- COMPANY: 	KOC UNIVERSITY
-- ENGINEER: 	ONURHAN OZTURK
-- 
-- CREATE DATE:    18:21:21 04/26/2016 
-- DESIGN NAME: 	
-- MODULE NAME:    SSSLIB - BEHAVIORAL 
-- PROJECT NAME: 	 SSSLIB
-- TARGET DEVICES: SPARTAN 3E
-- TOOL VERSIONS: 
-- DESCRIPTION: 
--		SSSLIB , Simple Seven Segment Library
--		is designed to add simple multiplexing 
--		solution to 4 digit seven segment displays.
--
-- DEPENDENCIES: 
--		SEVSEG_DRIVER.VHD
--		SEVSEG_DECODER.VHD
--		HUNDREDHZ_CLOCK_GENERATOR.VHD
--
-- REVISION:  A
-- REVISION 0.01 - FILE CREATED
-- ADDITIONAL COMMENTS: 
--		sozturk13@ku.edu.tr
--
----------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

-- UNCOMMENT THE FOLLOWING LIBRARY DECLARATION IF USING
-- ARITHMETIC FUNCTIONS WITH SIGNED OR UNSIGNED VALUES
--USE IEEE.NUMERIC_STD.ALL;

-- UNCOMMENT THE FOLLOWING LIBRARY DECLARATION IF INSTANTIATING
-- ANY XILINX PRIMITIVES IN THIS CODE.
--LIBRARY UNISIM;
--USE UNISIM.VCOMPONENTS.ALL;

ENTITY SSSLIB IS
    PORT ( A : IN  STD_LOGIC_VECTOR (4 DOWNTO 0);
           B : IN  STD_LOGIC_VECTOR (4 DOWNTO 0);
           C : IN  STD_LOGIC_VECTOR (4 DOWNTO 0);
           D : IN  STD_LOGIC_VECTOR (4 DOWNTO 0);
           MCLK : IN  STD_LOGIC;
           SEVSEG_DATA : OUT  STD_LOGIC_VECTOR (6 DOWNTO 0);
           SEVSEG_CONTROL : OUT  STD_LOGIC_VECTOR (7 DOWNTO 0));
END SSSLIB;

ARCHITECTURE BEHAVIORAL OF SSSLIB IS

--INTERMEDIATE SIGNALS
SIGNAL WIRE_HUNDREDHZ_CLOCK : STD_LOGIC;
SIGNAL WIRE_SEVSEG_DATA : STD_LOGIC_VECTOR(4 DOWNTO 0);

BEGIN

--ADD CLOCK GENERATOR
CLOCK_GENERATOR : ENTITY WORK.HUDREDHZ_CLOCK_GENERATOR PORT MAP(
	MCLK => MCLK,
	HUNDREDHZCLOCK => WIRE_HUNDREDHZ_CLOCK
);

--ADD DRIVER
DRIVER : ENTITY WORK.SEVSEG_DRIVER PORT MAP(
 A => A,
 B => B,
 C => C,
 D => D,
 CLK => WIRE_HUNDREDHZ_CLOCK,
 SEV_SEG_DATA => WIRE_SEVSEG_DATA,
 SEV_SEG_DRIVER => SEVSEG_CONTROL
);

--ADD DECODER
DECODER : ENTITY WORK.SEVSEG_DECODER PORT MAP(
	INPUT => WIRE_SEVSEG_DATA,
	SEVSEG_BUS => SEVSEG_DATA
);

END BEHAVIORAL;

